
`timescale 1ns/ 100ps
module b27s
	( (* altera_attribute = "-name IO_STANDARD \"3.3-V LVCMOS\"",    chip_pin = "49,46,25,24" *)
	input [3:0]sw,
	(* altera_attribute = "-name IO_STANDARD \"2.5V\"", useioff = 1, chip_pin = "67,68,69,70,71,72" *)
	output reg [6:0]led);
	
always @*
	case (sw)
		4'd0 : led = 7'b0111111;
		4'd1 : led = 7'b0000110;
		4'd2 : led = 7'b1011011;
		4'd3 : led = 7'b1001111;
		4'd4 : led = 7'b1100110;
		4'd5 : led = 7'b1101101;
		4'd6 : led = 7'b1111101;
		4'd7 : led = 7'b0000111;
		4'd8 : led = 7'b1111111;
		4'd9 : led = 7'b1101111;
		4'd10: led = 7'b1110111;
		4'd11: led = 7'b1111100;
		4'd12: led = 7'b0111001;
		4'd13: led = 7'b1011110;
		4'd14: led = 7'b1111011;
		4'd15: led = 7'b1110001;
	endcase
endmodule 	